entity test
end entity;